library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_pkg is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m.
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

(	7381	)	,
(	6320	)	,
(	6308	)	,
(	6296	)	,
(	6285	)	,
(	6273	)	,
(	6262	)	,
(	6250	)	,
(	6238	)	,
(	6227	)	, -- Element 9 of LUT
(	6215	)	,
(	6204	)	,
(	6192	)	,
(	6181	)	,
(	6169	)	,
(	6158	)	,
(	6147	)	,
(	6135	)	,
(	6124	)	,
(	6112	)	,
(	6101	)	, -- Element 20
(	6090	)	,
(	6078	)	,
(	6067	)	,
(	6056	)	,
(	6045	)	,
(	6033	)	,
(	6022	)	,
(	6011	)	,
(	6000	)	,
(	5989	)	,
(	5978	)	,
(	5967	)	,
(	5955	)	,
(	5944	)	,
(	5933	)	,
(	5922	)	,
(	5911	)	,
(	5900	)	,
(	5889	)	,
(	5878	)	,
(	5867	)	,
(	5856	)	,
(	5846	)	,
(	5835	)	,
(	5824	)	,
(	5813	)	,
(	5802	)	,
(	5791	)	,
(	5781	)	,
(	5770	)	,
(	5759	)	,
(	5748	)	,
(	5738	)	,
(	5727	)	,
(	5716	)	,
(	5706	)	,
(	5695	)	,
(	5684	)	,
(	5674	)	,
(	5663	)	,
(	5653	)	,
(	5642	)	,
(	5631	)	,
(	5621	)	,
(	5610	)	,
(	5600	)	,
(	5590	)	,
(	5579	)	,
(	5569	)	,
(	5558	)	,
(	5548	)	,
(	5537	)	,
(	5527	)	,
(	5517	)	,
(	5506	)	,
(	5496	)	,
(	5486	)	,
(	5476	)	,
(	5465	)	,
(	5455	)	,
(	5445	)	,
(	5435	)	,
(	5425	)	,
(	5414	)	,
(	5404	)	,
(	5394	)	,
(	5384	)	,
(	5374	)	,
(	5364	)	,
(	5354	)	,
(	5344	)	,
(	5334	)	,
(	5324	)	,
(	5314	)	,
(	5304	)	,
(	5294	)	,
(	5284	)	,
(	5274	)	,
(	5264	)	,
(	5254	)	,
(	5245	)	,
(	5235	)	,
(	5225	)	,
(	5215	)	,
(	5205	)	,
(	5195	)	,
(	5186	)	,
(	5176	)	,
(	5166	)	,
(	5157	)	,
(	5147	)	,
(	5137	)	,
(	5128	)	,
(	5118	)	,
(	5108	)	,
(	5099	)	,
(	5089	)	,
(	5080	)	,
(	5070	)	,
(	5061	)	,
(	5051	)	,
(	5042	)	,
(	5032	)	,
(	5023	)	,
(	5013	)	,
(	5004	)	,
(	4994	)	,
(	4985	)	,
(	4976	)	,
(	4966	)	,
(	4957	)	,
(	4947	)	,
(	4938	)	,
(	4929	)	,
(	4920	)	,
(	4910	)	,
(	4901	)	,
(	4892	)	,
(	4883	)	,
(	4873	)	,
(	4864	)	,
(	4855	)	,
(	4846	)	,
(	4837	)	,
(	4828	)	,
(	4819	)	,
(	4810	)	,
(	4800	)	,
(	4791	)	,
(	4782	)	,
(	4773	)	,
(	4764	)	,
(	4755	)	,
(	4746	)	,
(	4738	)	,
(	4729	)	,
(	4720	)	,
(	4711	)	,
(	4702	)	,
(	4693	)	,
(	4684	)	,
(	4675	)	,
(	4667	)	,
(	4658	)	,
(	4649	)	,
(	4640	)	,
(	4631	)	,
(	4623	)	,
(	4614	)	,
(	4605	)	,
(	4597	)	,
(	4588	)	,
(	4579	)	,
(	4571	)	,
(	4562	)	,
(	4553	)	,
(	4545	)	,
(	4536	)	,
(	4528	)	,
(	4519	)	,
(	4511	)	,
(	4502	)	,
(	4493	)	,
(	4485	)	,
(	4477	)	,
(	4468	)	,
(	4460	)	,
(	4451	)	,
(	4443	)	,
(	4434	)	,
(	4426	)	,
(	4418	)	,
(	4409	)	,
(	4401	)	,
(	4393	)	,
(	4384	)	,
(	4376	)	,
(	4368	)	,
(	4360	)	,
(	4351	)	,
(	4343	)	,
(	4335	)	,
(	4327	)	,
(	4319	)	,
(	4310	)	,
(	4302	)	,
(	4294	)	,
(	4286	)	,
(	4278	)	,
(	4270	)	,
(	4262	)	,
(	4254	)	,
(	4246	)	,
(	4238	)	,
(	4230	)	,
(	4222	)	,
(	4214	)	,
(	4206	)	,
(	4198	)	,
(	4190	)	,
(	4182	)	,
(	4174	)	,
(	4166	)	,
(	4158	)	,
(	4150	)	,
(	4142	)	,
(	4135	)	,
(	4127	)	,
(	4119	)	,
(	4111	)	,
(	4103	)	,
(	4096	)	,
(	4088	)	,
(	4080	)	,
(	4073	)	,
(	4065	)	,
(	4057	)	,
(	4049	)	,
(	4042	)	,
(	4034	)	,
(	4027	)	,
(	4019	)	,
(	4011	)	,
(	4004	)	,
(	3996	)	,
(	3989	)	,
(	3981	)	,
(	3974	)	,
(	3966	)	,
(	3959	)	,
(	3951	)	,
(	3944	)	,
(	3936	)	,
(	3929	)	,
(	3921	)	,
(	3914	)	,
(	3906	)	,
(	3899	)	,
(	3892	)	,
(	3884	)	,
(	3877	)	,
(	3870	)	,
(	3862	)	,
(	3855	)	,
(	3848	)	,
(	3841	)	,
(	3833	)	,
(	3826	)	,
(	3819	)	,
(	3812	)	,
(	3804	)	,
(	3797	)	,
(	3790	)	,
(	3783	)	,
(	3776	)	,
(	3769	)	,
(	3761	)	,
(	3754	)	,
(	3747	)	,
(	3740	)	,
(	3733	)	,
(	3726	)	,
(	3719	)	,
(	3712	)	,
(	3705	)	,
(	3698	)	,
(	3691	)	,
(	3684	)	,
(	3677	)	,
(	3670	)	,
(	3663	)	,
(	3656	)	,
(	3649	)	,
(	3643	)	,
(	3636	)	,
(	3629	)	,
(	3622	)	,
(	3615	)	,
(	3608	)	,
(	3602	)	,
(	3595	)	,
(	3588	)	,
(	3581	)	,
(	3574	)	,
(	3568	)	,
(	3561	)	,
(	3554	)	,
(	3548	)	,
(	3541	)	,
(	3534	)	,
(	3528	)	,
(	3521	)	,
(	3514	)	,
(	3508	)	,
(	3501	)	,
(	3494	)	,
(	3488	)	,
(	3481	)	,
(	3475	)	,
(	3468	)	,
(	3462	)	,
(	3455	)	,
(	3449	)	,
(	3442	)	,
(	3436	)	,
(	3429	)	,
(	3423	)	,
(	3416	)	,
(	3410	)	,
(	3404	)	,
(	3397	)	,
(	3391	)	,
(	3384	)	,
(	3378	)	,
(	3372	)	,
(	3365	)	,
(	3359	)	,
(	3353	)	,
(	3346	)	,
(	3340	)	,
(	3334	)	,
(	3328	)	,
(	3321	)	,
(	3315	)	,
(	3309	)	,
(	3303	)	,
(	3296	)	,
(	3290	)	,
(	3284	)	,
(	3278	)	,
(	3272	)	,
(	3266	)	,
(	3260	)	,
(	3253	)	,
(	3247	)	,
(	3241	)	,
(	3235	)	,
(	3229	)	,
(	3223	)	,
(	3217	)	,
(	3211	)	,
(	3205	)	,
(	3199	)	,
(	3193	)	,
(	3187	)	,
(	3181	)	,
(	3175	)	,
(	3169	)	,
(	3163	)	,
(	3157	)	,
(	3151	)	,
(	3146	)	,
(	3140	)	,
(	3134	)	,
(	3128	)	,
(	3122	)	,
(	3116	)	,
(	3110	)	,
(	3105	)	,
(	3099	)	,
(	3093	)	,
(	3087	)	,
(	3082	)	,
(	3076	)	,
(	3070	)	,
(	3064	)	,
(	3059	)	,
(	3053	)	,
(	3047	)	,
(	3042	)	,
(	3036	)	,
(	3030	)	,
(	3025	)	,
(	3019	)	,
(	3013	)	,
(	3008	)	,
(	3002	)	,
(	2997	)	,
(	2991	)	,
(	2985	)	,
(	2980	)	,
(	2974	)	,
(	2969	)	,
(	2963	)	,
(	2958	)	,
(	2952	)	,
(	2947	)	,
(	2941	)	,
(	2936	)	,
(	2931	)	,
(	2925	)	,
(	2920	)	,
(	2914	)	,
(	2909	)	,
(	2903	)	,
(	2898	)	,
(	2893	)	,
(	2887	)	,
(	2882	)	,
(	2877	)	,
(	2871	)	,
(	2866	)	,
(	2861	)	,
(	2855	)	,
(	2850	)	,
(	2845	)	,
(	2840	)	,
(	2834	)	,
(	2829	)	,
(	2824	)	,
(	2819	)	,
(	2814	)	,
(	2808	)	,
(	2803	)	,
(	2798	)	,
(	2793	)	,
(	2788	)	,
(	2783	)	,
(	2777	)	,
(	2772	)	,
(	2767	)	,
(	2762	)	,
(	2757	)	,
(	2752	)	,
(	2747	)	,
(	2742	)	,
(	2737	)	,
(	2732	)	,
(	2727	)	,
(	2722	)	,
(	2717	)	,
(	2712	)	,
(	2707	)	,
(	2702	)	,
(	2697	)	,
(	2692	)	,
(	2687	)	,
(	2682	)	,
(	2677	)	,
(	2672	)	,
(	2667	)	,
(	2663	)	,
(	2658	)	,
(	2653	)	,
(	2648	)	,
(	2643	)	,
(	2638	)	,
(	2634	)	,
(	2629	)	,
(	2624	)	,
(	2619	)	,
(	2614	)	,
(	2610	)	,
(	2605	)	,
(	2600	)	,
(	2595	)	,
(	2591	)	,
(	2586	)	,
(	2581	)	,
(	2577	)	,
(	2572	)	,
(	2567	)	,
(	2563	)	,
(	2558	)	,
(	2553	)	,
(	2549	)	,
(	2544	)	,
(	2539	)	,
(	2535	)	,
(	2530	)	,
(	2526	)	,
(	2521	)	,
(	2516	)	,
(	2512	)	,
(	2507	)	,
(	2503	)	,
(	2498	)	,
(	2494	)	,
(	2489	)	,
(	2485	)	,
(	2480	)	,
(	2476	)	,
(	2471	)	,
(	2467	)	,
(	2463	)	,
(	2458	)	,
(	2454	)	,
(	2449	)	,
(	2445	)	,
(	2440	)	,
(	2436	)	,
(	2432	)	,
(	2427	)	,
(	2423	)	,
(	2419	)	,
(	2414	)	,
(	2410	)	,
(	2406	)	,
(	2401	)	,
(	2397	)	,
(	2393	)	,
(	2388	)	,
(	2384	)	,
(	2380	)	,
(	2376	)	,
(	2371	)	,
(	2367	)	,
(	2363	)	,
(	2359	)	,
(	2355	)	,
(	2350	)	,
(	2346	)	,
(	2342	)	,
(	2338	)	,
(	2334	)	,
(	2330	)	,
(	2325	)	,
(	2321	)	,
(	2317	)	,
(	2313	)	,
(	2309	)	,
(	2305	)	,
(	2301	)	,
(	2297	)	,
(	2293	)	,
(	2289	)	,
(	2285	)	,
(	2281	)	,
(	2277	)	,
(	2272	)	,
(	2268	)	,
(	2264	)	,
(	2260	)	,
(	2257	)	,
(	2253	)	,
(	2249	)	,
(	2245	)	,
(	2241	)	,
(	2237	)	,
(	2233	)	,
(	2229	)	,
(	2225	)	,
(	2221	)	,
(	2217	)	,
(	2213	)	,
(	2209	)	,
(	2206	)	,
(	2202	)	,
(	2198	)	,
(	2194	)	,
(	2190	)	,
(	2186	)	,
(	2183	)	,
(	2179	)	,
(	2175	)	,
(	2171	)	,
(	2167	)	,
(	2164	)	,
(	2160	)	,
(	2156	)	,
(	2152	)	,
(	2149	)	,
(	2145	)	,
(	2141	)	,
(	2137	)	,
(	2134	)	,
(	2130	)	,
(	2126	)	,
(	2123	)	,
(	2119	)	,
(	2115	)	,
(	2112	)	,
(	2108	)	,
(	2104	)	,
(	2101	)	,
(	2097	)	,
(	2094	)	,
(	2090	)	,
(	2086	)	,
(	2083	)	,
(	2079	)	,
(	2076	)	,
(	2072	)	,
(	2069	)	,
(	2065	)	,
(	2061	)	,
(	2058	)	,
(	2054	)	,
(	2051	)	,
(	2047	)	,
(	2044	)	,
(	2040	)	,
(	2037	)	,
(	2033	)	,
(	2030	)	,
(	2027	)	,
(	2023	)	,
(	2020	)	,
(	2016	)	,
(	2013	)	,
(	2009	)	,
(	2006	)	,
(	2003	)	,
(	1999	)	,
(	1996	)	,
(	1992	)	,
(	1989	)	,
(	1986	)	,
(	1982	)	,
(	1979	)	,
(	1976	)	,
(	1972	)	,
(	1969	)	,
(	1966	)	,
(	1962	)	,
(	1959	)	,
(	1956	)	,
(	1953	)	,
(	1949	)	,
(	1946	)	,
(	1943	)	,
(	1940	)	,
(	1936	)	,
(	1933	)	,
(	1930	)	,
(	1927	)	,
(	1923	)	,
(	1920	)	,
(	1917	)	,
(	1914	)	,
(	1911	)	,
(	1907	)	,
(	1904	)	,
(	1901	)	,
(	1898	)	,
(	1895	)	,
(	1892	)	,
(	1889	)	,
(	1885	)	,
(	1882	)	,
(	1879	)	,
(	1876	)	,
(	1873	)	,
(	1870	)	,
(	1867	)	,
(	1864	)	,
(	1861	)	,
(	1858	)	,
(	1855	)	,
(	1852	)	,
(	1849	)	,
(	1846	)	,
(	1843	)	,
(	1840	)	,
(	1836	)	,
(	1834	)	,
(	1831	)	,
(	1828	)	,
(	1825	)	,
(	1822	)	,
(	1819	)	,
(	1816	)	,
(	1813	)	,
(	1810	)	,
(	1807	)	,
(	1804	)	,
(	1801	)	,
(	1798	)	,
(	1795	)	,
(	1792	)	,
(	1789	)	,
(	1787	)	,
(	1784	)	,
(	1781	)	,
(	1778	)	,
(	1775	)	,
(	1772	)	,
(	1769	)	,
(	1767	)	,
(	1764	)	,
(	1761	)	,
(	1758	)	,
(	1755	)	,
(	1752	)	,
(	1750	)	,
(	1747	)	,
(	1744	)	,
(	1741	)	,
(	1739	)	,
(	1736	)	,
(	1733	)	,
(	1730	)	,
(	1728	)	,
(	1725	)	,
(	1722	)	,
(	1719	)	,
(	1717	)	,
(	1714	)	,
(	1711	)	,
(	1709	)	,
(	1706	)	,
(	1703	)	,
(	1701	)	,
(	1698	)	,
(	1695	)	,
(	1693	)	,
(	1690	)	,
(	1687	)	,
(	1685	)	,
(	1682	)	,
(	1679	)	,
(	1677	)	,
(	1674	)	,
(	1672	)	,
(	1669	)	,
(	1666	)	,
(	1664	)	,
(	1661	)	,
(	1659	)	,
(	1656	)	,
(	1654	)	,
(	1651	)	,
(	1648	)	,
(	1646	)	,
(	1643	)	,
(	1641	)	,
(	1638	)	,
(	1636	)	,
(	1633	)	,
(	1631	)	,
(	1628	)	,
(	1626	)	,
(	1623	)	,
(	1621	)	,
(	1618	)	,
(	1616	)	,
(	1613	)	,
(	1611	)	,
(	1609	)	,
(	1606	)	,
(	1604	)	,
(	1601	)	,
(	1599	)	,
(	1596	)	,
(	1594	)	,
(	1592	)	,
(	1589	)	,
(	1587	)	,
(	1584	)	,
(	1582	)	,
(	1580	)	,
(	1577	)	,
(	1575	)	,
(	1573	)	,
(	1570	)	,
(	1568	)	,
(	1566	)	,
(	1563	)	,
(	1561	)	,
(	1559	)	,
(	1556	)	,
(	1554	)	,
(	1552	)	,
(	1549	)	,
(	1547	)	,
(	1545	)	,
(	1543	)	,
(	1540	)	,
(	1538	)	,
(	1536	)	,
(	1533	)	,
(	1531	)	,
(	1529	)	,
(	1527	)	,
(	1525	)	,
(	1522	)	,
(	1520	)	,
(	1518	)	,
(	1516	)	,
(	1513	)	,
(	1511	)	,
(	1509	)	,
(	1507	)	,
(	1505	)	,
(	1502	)	,
(	1500	)	,
(	1498	)	,
(	1496	)	,
(	1494	)	,
(	1492	)	,
(	1490	)	,
(	1487	)	,
(	1485	)	,
(	1483	)	,
(	1481	)	,
(	1479	)	,
(	1477	)	,
(	1475	)	,
(	1473	)	,
(	1470	)	,
(	1468	)	,
(	1466	)	,
(	1464	)	,
(	1462	)	,
(	1460	)	,
(	1458	)	,
(	1456	)	,
(	1454	)	,
(	1452	)	,
(	1450	)	,
(	1448	)	,
(	1446	)	,
(	1444	)	,
(	1442	)	,
(	1440	)	,
(	1438	)	,
(	1436	)	,
(	1434	)	,
(	1432	)	,
(	1430	)	,
(	1428	)	,
(	1426	)	,
(	1424	)	,
(	1422	)	,
(	1420	)	,
(	1418	)	,
(	1416	)	,
(	1414	)	,
(	1412	)	,
(	1410	)	,
(	1408	)	,
(	1406	)	,
(	1404	)	,
(	1402	)	,
(	1400	)	,
(	1398	)	,
(	1397	)	,
(	1395	)	,
(	1393	)	,
(	1391	)	,
(	1389	)	,
(	1387	)	,
(	1385	)	,
(	1383	)	,
(	1381	)	,
(	1380	)	,
(	1378	)	,
(	1376	)	,
(	1374	)	,
(	1372	)	,
(	1370	)	,
(	1368	)	,
(	1367	)	,
(	1365	)	,
(	1363	)	,
(	1361	)	,
(	1359	)	,
(	1358	)	,
(	1356	)	,
(	1354	)	,
(	1352	)	,
(	1350	)	,
(	1349	)	,
(	1347	)	,
(	1345	)	,
(	1343	)	,
(	1342	)	,
(	1340	)	,
(	1338	)	,
(	1336	)	,
(	1335	)	,
(	1333	)	,
(	1331	)	,
(	1329	)	,
(	1328	)	,
(	1326	)	,
(	1324	)	,
(	1322	)	,
(	1321	)	,
(	1319	)	,
(	1317	)	,
(	1316	)	,
(	1314	)	,
(	1312	)	,
(	1311	)	,
(	1309	)	,
(	1307	)	,
(	1305	)	,
(	1304	)	,
(	1302	)	,
(	1300	)	,
(	1299	)	,
(	1297	)	,
(	1296	)	,
(	1294	)	,
(	1292	)	,
(	1291	)	,
(	1289	)	,
(	1287	)	,
(	1286	)	,
(	1284	)	,
(	1283	)	,
(	1281	)	,
(	1279	)	,
(	1278	)	,
(	1276	)	,
(	1275	)	,
(	1273	)	,
(	1271	)	,
(	1270	)	,
(	1268	)	,
(	1267	)	,
(	1265	)	,
(	1264	)	,
(	1262	)	,
(	1260	)	,
(	1259	)	,
(	1257	)	,
(	1256	)	,
(	1254	)	,
(	1253	)	,
(	1251	)	,
(	1250	)	,
(	1248	)	,
(	1247	)	,
(	1245	)	,
(	1244	)	,
(	1242	)	,
(	1241	)	,
(	1239	)	,
(	1238	)	,
(	1236	)	,
(	1235	)	,
(	1233	)	,
(	1232	)	,
(	1230	)	,
(	1229	)	,
(	1227	)	,
(	1226	)	,
(	1224	)	,
(	1223	)	,
(	1221	)	,
(	1220	)	,
(	1218	)	,
(	1217	)	,
(	1216	)	,
(	1214	)	,
(	1213	)	,
(	1211	)	,
(	1210	)	,
(	1208	)	,
(	1207	)	,
(	1206	)	,
(	1204	)	,
(	1203	)	,
(	1201	)	,
(	1200	)	,
(	1199	)	,
(	1197	)	,
(	1196	)	,
(	1194	)	,
(	1193	)	,
(	1192	)	,
(	1190	)	,
(	1189	)	,
(	1188	)	,
(	1186	)	,
(	1185	)	,
(	1184	)	,
(	1182	)	,
(	1181	)	,
(	1179	)	,
(	1178	)	,
(	1177	)	,
(	1175	)	,
(	1174	)	,
(	1173	)	,
(	1171	)	,
(	1170	)	,
(	1169	)	,
(	1168	)	,
(	1166	)	,
(	1165	)	,
(	1164	)	,
(	1162	)	,
(	1161	)	,
(	1160	)	,
(	1158	)	,
(	1157	)	,
(	1156	)	,
(	1155	)	,
(	1153	)	,
(	1152	)	,
(	1151	)	,
(	1149	)	,
(	1148	)	,
(	1147	)	,
(	1146	)	,
(	1144	)	,
(	1143	)	,
(	1142	)	,
(	1141	)	,
(	1139	)	,
(	1138	)	,
(	1137	)	,
(	1136	)	,
(	1135	)	,
(	1133	)	,
(	1132	)	,
(	1131	)	,
(	1130	)	,
(	1128	)	,
(	1127	)	,
(	1126	)	,
(	1125	)	,
(	1124	)	,
(	1122	)	,
(	1121	)	,
(	1120	)	,
(	1119	)	,
(	1118	)	,
(	1116	)	,
(	1115	)	,
(	1114	)	,
(	1113	)	,
(	1112	)	,
(	1111	)	,
(	1109	)	,
(	1108	)	,
(	1107	)	,
(	1106	)	,
(	1105	)	,
(	1104	)	,
(	1103	)	,
(	1101	)	,
(	1100	)	,
(	1099	)	,
(	1098	)	,
(	1097	)	,
(	1096	)	,
(	1095	)	,
(	1093	)	,
(	1092	)	,
(	1091	)	,
(	1090	)	,
(	1089	)	,
(	1088	)	,
(	1087	)	,
(	1086	)	,
(	1085	)	,
(	1083	)	,
(	1082	)	,
(	1081	)	,
(	1080	)	,
(	1079	)	,
(	1078	)	,
(	1077	)	,
(	1076	)	,
(	1075	)	,
(	1074	)	,
(	1073	)	,
(	1072	)	,
(	1070	)	,
(	1069	)	,
(	1068	)	,
(	1067	)	,
(	1066	)	,
(	1065	)	,
(	1064	)	,
(	1063	)	,
(	1062	)	,
(	1061	)	,
(	1060	)	,
(	1059	)	,
(	1058	)	,
(	1057	)	,
(	1056	)	,
(	1055	)	,
(	1054	)	,
(	1053	)	,
(	1052	)	,
(	1051	)	,
(	1050	)	,
(	1049	)	,
(	1048	)	,
(	1047	)	,
(	1046	)	,
(	1045	)	,
(	1044	)	,
(	1043	)	,
(	1042	)	,
(	1041	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1037	)	,
(	1036	)	,
(	1035	)	,
(	1034	)	,
(	1033	)	,
(	1032	)	,
(	1031	)	,
(	1030	)	,
(	1029	)	,
(	1028	)	,
(	1027	)	,
(	1026	)	,
(	1025	)	,
(	1024	)	,
(	1023	)	,
(	1022	)	,
(	1021	)	,
(	1020	)	,
(	1019	)	,
(	1018	)	,
(	1018	)	,
(	1017	)	,
(	1016	)	,
(	1015	)	,
(	1014	)	,
(	1013	)	,
(	1012	)	,
(	1011	)	,
(	1010	)	,
(	1009	)	,
(	1008	)	,
(	1007	)	,
(	1006	)	,
(	1006	)	,
(	1005	)	,
(	1004	)	,
(	1003	)	,
(	1002	)	,
(	1001	)	,
(	1000	)	,
(	999	)	,
(	998	)	,
(	997	)	,
(	997	)	,
(	996	)	,
(	995	)	,
(	994	)	,
(	993	)	,
(	992	)	,
(	991	)	,
(	990	)	,
(	990	)	,
(	989	)	,
(	988	)	,
(	987	)	,
(	986	)	,
(	985	)	,
(	984	)	,
(	983	)	,
(	983	)	,
(	982	)	,
(	981	)	,
(	980	)	,
(	979	)	,
(	978	)	,
(	977	)	,
(	977	)	,
(	976	)	,
(	975	)	,
(	974	)	,
(	973	)	,
(	972	)	,
(	972	)	,
(	971	)	,
(	970	)	,
(	969	)	,
(	968	)	,
(	967	)	,
(	967	)	,
(	966	)	,
(	965	)	,
(	964	)	,
(	963	)	,
(	963	)	,
(	962	)	,
(	961	)	,
(	960	)	,
(	959	)	,
(	959	)	,
(	958	)	,
(	957	)	,
(	956	)	,
(	955	)	,
(	955	)	,
(	954	)	,
(	953	)	,
(	952	)	,
(	951	)	,
(	951	)	,
(	950	)	,
(	949	)	,
(	948	)	,
(	947	)	,
(	947	)	,
(	946	)	,
(	945	)	,
(	944	)	,
(	944	)	,
(	943	)	,
(	942	)	,
(	941	)	,
(	941	)	,
(	940	)	,
(	939	)	,
(	938	)	,
(	937	)	,
(	937	)	,
(	936	)	,
(	935	)	,
(	934	)	,
(	934	)	,
(	933	)	,
(	932	)	,
(	931	)	,
(	931	)	,
(	930	)	,
(	929	)	,
(	928	)	,
(	928	)	,
(	927	)	,
(	926	)	,
(	925	)	,
(	925	)	,
(	924	)	,
(	923	)	,
(	923	)	,
(	922	)	,
(	921	)	,
(	920	)	,
(	920	)	,
(	919	)	,
(	918	)	,
(	917	)	,
(	917	)	,
(	916	)	,
(	915	)	,
(	915	)	,
(	914	)	,
(	913	)	,
(	912	)	,
(	912	)	,
(	911	)	,
(	910	)	,
(	910	)	,
(	909	)	,
(	908	)	,
(	908	)	,
(	907	)	,
(	906	)	,
(	905	)	,
(	905	)	,
(	904	)	,
(	903	)	,
(	903	)	,
(	902	)	,
(	901	)	,
(	901	)	,
(	900	)	,
(	899	)	,
(	899	)	,
(	898	)	,
(	897	)	,
(	896	)	,
(	896	)	,
(	895	)	,
(	894	)	,
(	894	)	,
(	893	)	,
(	892	)	,
(	892	)	,
(	891	)	,
(	890	)	,
(	890	)	,
(	889	)	,
(	888	)	,
(	888	)	,
(	887	)	,
(	886	)	,
(	886	)	,
(	885	)	,
(	884	)	,
(	884	)	,
(	883	)	,
(	882	)	,
(	882	)	,
(	881	)	,
(	880	)	,
(	880	)	,
(	879	)	,
(	878	)	,
(	878	)	,
(	877	)	,
(	877	)	,
(	876	)	,
(	875	)	,
(	875	)	,
(	874	)	,
(	873	)	,
(	873	)	,
(	872	)	,
(	871	)	,
(	871	)	,
(	870	)	,
(	869	)	,
(	869	)	,
(	868	)	,
(	868	)	,
(	867	)	,
(	866	)	,
(	866	)	,
(	865	)	,
(	864	)	,
(	864	)	,
(	863	)	,
(	862	)	,
(	862	)	,
(	861	)	,
(	861	)	,
(	860	)	,
(	859	)	,
(	859	)	,
(	858	)	,
(	857	)	,
(	857	)	,
(	856	)	,
(	856	)	,
(	855	)	,
(	854	)	,
(	854	)	,
(	853	)	,
(	853	)	,
(	852	)	,
(	851	)	,
(	851	)	,
(	850	)	,
(	849	)	,
(	849	)	,
(	848	)	,
(	848	)	,
(	847	)	,
(	846	)	,
(	846	)	,
(	845	)	,
(	845	)	,
(	844	)	,
(	843	)	,
(	843	)	,
(	842	)	,
(	842	)	,
(	841	)	,
(	840	)	,
(	840	)	,
(	839	)	,
(	839	)	,
(	838	)	,
(	837	)	,
(	837	)	,
(	836	)	,
(	836	)	,
(	835	)	,
(	834	)	,
(	834	)	,
(	833	)	,
(	833	)	,
(	832	)	,
(	832	)	,
(	831	)	,
(	830	)	,
(	830	)	,
(	829	)	,
(	829	)	,
(	828	)	,
(	827	)	,
(	827	)	,
(	826	)	,
(	826	)	,
(	825	)	,
(	824	)	,
(	824	)	,
(	823	)	,
(	823	)	,
(	822	)	,
(	822	)	,
(	821	)	,
(	820	)	,
(	820	)	,
(	819	)	,
(	819	)	,
(	818	)	,
(	818	)	,
(	817	)	,
(	816	)	,
(	816	)	,
(	815	)	,
(	815	)	,
(	814	)	,
(	814	)	,
(	813	)	,
(	812	)	,
(	812	)	,
(	811	)	,
(	811	)	,
(	810	)	,
(	810	)	,
(	809	)	,
(	808	)	,
(	808	)	,
(	807	)	,
(	807	)	,
(	806	)	,
(	806	)	,
(	805	)	,
(	805	)	,
(	804	)	,
(	803	)	,
(	803	)	,
(	802	)	,
(	802	)	,
(	801	)	,
(	801	)	,
(	800	)	,
(	799	)	,
(	799	)	,
(	798	)	,
(	798	)	,
(	797	)	,
(	797	)	,
(	796	)	,
(	796	)	,
(	795	)	,
(	794	)	,
(	794	)	,
(	793	)	,
(	793	)	,
(	792	)	,
(	792	)	,
(	791	)	,
(	791	)	,
(	790	)	,
(	790	)	,
(	789	)	,
(	788	)	,
(	788	)	,
(	787	)	,
(	787	)	,
(	786	)	,
(	786	)	,
(	785	)	,
(	785	)	,
(	784	)	,
(	784	)	,
(	783	)	,
(	782	)	,
(	782	)	,
(	781	)	,
(	781	)	,
(	780	)	,
(	780	)	,
(	779	)	,
(	779	)	,
(	778	)	,
(	778	)	,
(	777	)	,
(	776	)	,
(	776	)	,
(	775	)	,
(	775	)	,
(	774	)	,
(	774	)	,
(	773	)	,
(	773	)	,
(	772	)	,
(	772	)	,
(	771	)	,
(	770	)	,
(	770	)	,
(	769	)	,
(	769	)	,
(	768	)	,
(	768	)	,
(	767	)	,
(	767	)	,
(	766	)	,
(	766	)	,
(	765	)	,
(	765	)	,
(	764	)	,
(	764	)	,
(	763	)	,
(	762	)	,
(	762	)	,
(	761	)	,
(	761	)	,
(	760	)	,
(	760	)	,
(	759	)	,
(	759	)	,
(	758	)	,
(	758	)	,
(	757	)	,
(	757	)	,
(	756	)	,
(	756	)	,
(	755	)	,
(	754	)	,
(	754	)	,
(	753	)	,
(	753	)	,
(	752	)	,
(	752	)	,
(	751	)	,
(	751	)	,
(	750	)	,
(	750	)	,
(	749	)	,
(	749	)	,
(	748	)	,
(	748	)	,
(	747	)	,
(	746	)	,
(	746	)	,
(	745	)	,
(	745	)	,
(	744	)	,
(	744	)	,
(	743	)	,
(	743	)	,
(	742	)	,
(	742	)	,
(	741	)	,
(	741	)	,
(	740	)	,
(	740	)	,
(	739	)	,
(	739	)	,
(	738	)	,
(	737	)	,
(	737	)	,
(	736	)	,
(	736	)	,
(	735	)	,
(	735	)	,
(	734	)	,
(	734	)	,
(	733	)	,
(	733	)	,
(	732	)	,
(	732	)	,
(	731	)	,
(	731	)	,
(	730	)	,
(	730	)	,
(	729	)	,
(	729	)	,
(	728	)	,
(	727	)	,
(	727	)	,
(	726	)	,
(	726	)	,
(	725	)	,
(	725	)	,
(	724	)	,
(	724	)	,
(	723	)	,
(	723	)	,
(	722	)	,
(	722	)	,
(	721	)	,
(	721	)	,
(	720	)	,
(	720	)	,
(	719	)	,
(	719	)	,
(	718	)	,
(	718	)	,
(	717	)	,
(	716	)	,
(	716	)	,
(	715	)	,
(	715	)	,
(	714	)	,
(	714	)	,
(	713	)	,
(	713	)	,
(	712	)	,
(	712	)	,
(	711	)	,
(	711	)	,
(	710	)	,
(	710	)	,
(	709	)	,
(	709	)	,
(	708	)	,
(	708	)	,
(	707	)	,
(	707	)	,
(	706	)	,
(	705	)	,
(	705	)	,
(	704	)	,
(	704	)	,
(	703	)	,
(	703	)	,
(	702	)	,
(	702	)	,
(	701	)	,
(	701	)	,
(	700	)	,
(	700	)	,
(	699	)	,
(	699	)	,
(	698	)	,
(	698	)	,
(	697	)	,
(	697	)	,
(	696	)	,
(	696	)	,
(	695	)	,
(	694	)	,
(	694	)	,
(	693	)	,
(	693	)	,
(	692	)	,
(	692	)	,
(	691	)	,
(	691	)	,
(	690	)	,
(	690	)	,
(	689	)	,
(	689	)	,
(	688	)	,
(	688	)	,
(	687	)	,
(	687	)	,
(	686	)	,
(	686	)	,
(	685	)	,
(	685	)	,
(	684	)	,
(	683	)	,
(	683	)	,
(	682	)	,
(	682	)	,
(	681	)	,
(	681	)	,
(	680	)	,
(	680	)	,
(	679	)	,
(	679	)	,
(	678	)	,
(	678	)	,
(	677	)	,
(	677	)	,
(	676	)	,
(	676	)	,
(	675	)	,
(	675	)	,
(	674	)	,
(	673	)	,
(	673	)	,
(	672	)	,
(	672	)	,
(	671	)	,
(	671	)	,
(	670	)	,
(	670	)	,
(	669	)	,
(	669	)	,
(	668	)	,
(	668	)	,
(	667	)	,
(	667	)	,
(	666	)	,
(	666	)	,
(	665	)	,
(	665	)	,
(	664	)	,
(	663	)	,
(	663	)	,
(	662	)	,
(	662	)	,
(	661	)	,
(	661	)	,
(	660	)	,
(	660	)	,
(	659	)	,
(	659	)	,
(	658	)	,
(	658	)	,
(	657	)	,
(	657	)	,
(	656	)	,
(	656	)	,
(	655	)	,
(	655	)	,
(	654	)	,
(	653	)	,
(	653	)	,
(	652	)	,
(	652	)	,
(	651	)	,
(	651	)	,
(	650	)	,
(	650	)	,
(	649	)	,
(	649	)	,
(	648	)	,
(	648	)	,
(	647	)	,
(	647	)	,
(	646	)	,
(	646	)	,
(	645	)	,
(	645	)	,
(	644	)	,
(	643	)	,
(	643	)	,
(	642	)	,
(	642	)	,
(	641	)	,
(	641	)	,
(	640	)	,
(	640	)	,
(	639	)	,
(	639	)	,
(	638	)	,
(	638	)	,
(	637	)	,
(	637	)	,
(	636	)	,
(	636	)	,
(	635	)	,
(	634	)	,
(	634	)	,
(	633	)	,
(	633	)	,
(	632	)	,
(	632	)	,
(	631	)	,
(	631	)	,
(	630	)	,
(	630	)	,
(	629	)	,
(	629	)	,
(	628	)	,
(	628	)	,
(	627	)	,
(	627	)	,
(	626	)	,
(	625	)	,
(	625	)	,
(	624	)	,
(	624	)	,
(	623	)	,
(	623	)	,
(	622	)	,
(	622	)	,
(	621	)	,
(	621	)	,
(	620	)	,
(	620	)	,
(	619	)	,
(	619	)	,
(	618	)	,
(	618	)	,
(	617	)	,
(	616	)	,
(	616	)	,
(	615	)	,
(	615	)	,
(	614	)	,
(	614	)	,
(	613	)	,
(	613	)	,
(	612	)	,
(	612	)	,
(	611	)	,
(	611	)	,
(	610	)	,
(	610	)	,
(	609	)	,
(	608	)	,
(	608	)	,
(	607	)	,
(	607	)	,
(	606	)	,
(	606	)	,
(	605	)	,
(	605	)	,
(	604	)	,
(	604	)	,
(	603	)	,
(	603	)	,
(	602	)	,
(	602	)	,
(	601	)	,
(	601	)	,
(	600	)	,
(	599	)	,
(	599	)	,
(	598	)	,
(	598	)	,
(	597	)	,
(	597	)	,
(	596	)	,
(	596	)	,
(	595	)	,
(	595	)	,
(	594	)	,
(	594	)	,
(	593	)	,
(	593	)	,
(	592	)	,
(	592	)	,
(	591	)	,
(	590	)	,
(	590	)	,
(	589	)	,
(	589	)	,
(	588	)	,
(	588	)	,
(	587	)	,
(	587	)	,
(	586	)	,
(	586	)	,
(	585	)	,
(	585	)	,
(	584	)	,
(	584	)	,
(	583	)	,
(	583	)	,
(	582	)	,
(	581	)	,
(	581	)	,
(	580	)	,
(	580	)	,
(	579	)	,
(	579	)	,
(	578	)	,
(	578	)	,
(	577	)	,
(	577	)	,
(	576	)	,
(	576	)	,
(	575	)	,
(	575	)	,
(	574	)	,
(	574	)	,
(	573	)	,
(	572	)	,
(	572	)	,
(	571	)	,
(	571	)	,
(	570	)	,
(	570	)	,
(	569	)	,
(	569	)	,
(	568	)	,
(	568	)	,
(	567	)	,
(	567	)	,
(	566	)	,
(	566	)	,
(	565	)	,
(	565	)	,
(	564	)	,
(	564	)	,
(	563	)	,
(	562	)	,
(	562	)	,
(	561	)	,
(	561	)	,
(	560	)	,
(	560	)	,
(	559	)	,
(	559	)	,
(	558	)	,
(	558	)	,
(	557	)	,
(	557	)	,
(	556	)	,
(	556	)	,
(	555	)	,
(	555	)	,
(	554	)	,
(	554	)	,
(	553	)	,
(	553	)	,
(	552	)	,
(	551	)	,
(	551	)	,
(	550	)	,
(	550	)	,
(	549	)	,
(	549	)	,
(	548	)	,
(	548	)	,
(	547	)	,
(	547	)	,
(	546	)	,
(	546	)	,
(	545	)	,
(	545	)	,
(	544	)	,
(	544	)	,
(	543	)	,
(	543	)	,
(	542	)	,
(	542	)	,
(	541	)	,
(	541	)	,
(	540	)	,
(	540	)	,
(	539	)	,
(	538	)	,
(	538	)	,
(	537	)	,
(	537	)	,
(	536	)	,
(	536	)	,
(	535	)	,
(	535	)	,
(	534	)	,
(	534	)	,
(	533	)	,
(	533	)	,
(	532	)	,
(	532	)	,
(	531	)	,
(	531	)	,
(	530	)	,
(	530	)	,
(	529	)	,
(	529	)	,
(	528	)	,
(	528	)	,
(	527	)	,
(	527	)	,
(	526	)	,
(	526	)	,
(	525	)	,
(	525	)	,
(	524	)	,
(	524	)	,
(	523	)	,
(	523	)	,
(	522	)	,
(	522	)	,
(	521	)	,
(	521	)	,
(	520	)	,
(	520	)	,
(	519	)	,
(	519	)	,
(	518	)	,
(	518	)	,
(	517	)	,
(	517	)	,
(	516	)	,
(	516	)	,
(	515	)	,
(	515	)	,
(	514	)	,
(	514	)	,
(	513	)	,
(	513	)	,
(	512	)	,
(	512	)	,
(	511	)	,
(	511	)	,
(	510	)	,
(	510	)	,
(	509	)	,
(	509	)	,
(	508	)	,
(	508	)	,
(	507	)	,
(	507	)	,
(	506	)	,
(	506	)	,
(	505	)	,
(	505	)	,
(	504	)	,
(	504	)	,
(	503	)	,
(	503	)	,
(	502	)	,
(	502	)	,
(	501	)	,
(	501	)	,
(	500	)	,
(	500	)	,
(	499	)	,
(	499	)	,
(	498	)	,
(	498	)	,
(	497	)	,
(	497	)	,
(	496	)	,
(	496	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	494	)	,
(	494	)	,
(	493	)	,
(	493	)	,
(	492	)	,
(	492	)	,
(	491	)	,
(	491	)	,
(	490	)	,
(	490	)	,
(	489	)	,
(	489	)	,
(	488	)	,
(	488	)	,
(	487	)	,
(	487	)	,
(	486	)	,
(	486	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	484	)	,
(	484	)	,
(	483	)	,
(	483	)	,
(	482	)	,
(	482	)	,
(	481	)	,
(	481	)	,
(	480	)	,
(	480	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	478	)	,
(	478	)	,
(	477	)	,
(	477	)	,
(	476	)	,
(	476	)	,
(	475	)	,
(	475	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	473	)	,
(	473	)	,
(	472	)	,
(	472	)	,
(	471	)	,
(	471	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	469	)	,
(	469	)	,
(	468	)	,
(	468	)	,
(	467	)	,
(	467	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	465	)	,
(	465	)	,
(	464	)	,
(	464	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	462	)	,
(	462	)	,
(	461	)	,
(	461	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	459	)	,
(	459	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	457	)	,
(	457	)	,
(	456	)	,
(	456	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	454	)	,
(	454	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	452	)	,
(	452	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	450	)	,
(	450	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	448	)	,
(	448	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	446	)	,
(	446	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	443	)	,
(	443	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	441	)	,
(	441	)	,
(	441	)	,
(	440	)	,
(	440	)	,
(	439	)	,
(	439	)	,
(	439	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	436	)	,
(	436	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	433	)	,
(	433	)	,
(	433	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	429	)	,
(	429	)	,
(	429	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	425	)	,
(	425	)	,
(	425	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	419	)	,
(	419	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	422	)	,
(	422	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	424	)	,
(	424	)	,
(	425	)	,
(	425	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	427	)	,
(	427	)	,
(	428	)	,
(	428	)	,
(	429	)	,
(	429	)	,
(	430	)	,
(	430	)	,
(	431	)	,
(	431	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	433	)	,
(	433	)	,
(	434	)	,
(	434	)	,
(	435	)	,
(	435	)	,
(	436	)	,
(	437	)	,
(	437	)	,
(	438	)	,
(	438	)	,
(	439	)	,
(	439	)	,
(	440	)	,
(	440	)	,
(	441	)	,
(	441	)	,
(	442	)	,
(	443	)	,
(	443	)	,
(	444	)	,
(	444	)	,
(	445	)	,
(	445	)	,
(	446	)	,
(	447	)	,
(	447	)	,
(	448	)	,
(	448	)	,
(	449	)	,
(	450	)	,
(	450	)	,
(	451	)	,
(	451	)	,
(	452	)	,
(	453	)	,
(	453	)	,
(	454	)	,
(	455	)	,
(	455	)	,
(	456	)	,
(	457	)	,
(	457	)	,
(	458	)	,
(	459	)	,
(	459	)	,
(	460	)	,
(	461	)	,
(	461	)	,
(	462	)	,
(	463	)	,
(	464	)	,
(	464	)	,
(	465	)	,
(	466	)	,
(	466	)	,
(	467	)	,
(	468	)	,
(	469	)	,
(	469	)	,
(	470	)	,
(	471	)	,
(	472	)	,
(	472	)	,
(	473	)	,
(	474	)	,
(	475	)	,
(	476	)	,
(	476	)	,
(	477	)	,
(	478	)	,
(	479	)	,
(	480	)	,
(	480	)	,
(	481	)	,
(	482	)	,
(	483	)	,
(	484	)	,
(	485	)	,
(	485	)	,
(	486	)	,
(	487	)	,
(	488	)	,
(	489	)	,
(	490	)	,
(	491	)	,
(	491	)	,
(	492	)	,
(	493	)	,
(	494	)	,
(	495	)	,
(	496	)	,
(	497	)	,
(	498	)	,
(	499	)	,
(	500	)	,
(	500	)	,
(	501	)	,
(	502	)	,
(	503	)	,
(	504	)	,
(	505	)	,
(	506	)	,
(	507	)	,
(	508	)	,
(	509	)	,
(	510	)	,
(	511	)	,
(	512	)	,
(	513	)	,
(	514	)	,
(	515	)	,
(	516	)	,
(	517	)	,
(	518	)	,
(	519	)	,
(	520	)	,
(	521	)	,
(	522	)	,
(	523	)	,
(	524	)	,
(	525	)	,
(	526	)	,
(	527	)	,
(	528	)	,
(	530	)	,
(	531	)	,
(	532	)	,
(	533	)	,
(	534	)	,
(	535	)	,
(	536	)	,
(	537	)	,
(	538	)	,
(	540	)	,
(	541	)	,
(	542	)	,
(	543	)	,
(	544	)	,
(	545	)	,
(	546	)	,
(	548	)	,
(	549	)	,
(	550	)	,
(	551	)	,
(	552	)	,
(	553	)	,
(	555	)	,
(	556	)	,
(	557	)	,
(	558	)	,
(	560	)	,
(	561	)	,
(	562	)	,
(	563	)	,
(	565	)	,
(	566	)	,
(	567	)	,
(	568	)	,
(	570	)	,
(	571	)	,
(	572	)	,
(	573	)	,
(	575	)	,
(	576	)	,
(	577	)	,
(	579	)	,
(	580	)	,
(	581	)	,
(	583	)	,
(	584	)	,
(	585	)	,
(	587	)	,
(	588	)	,
(	589	)	,
(	591	)	,
(	592	)	,
(	593	)	,
(	595	)	,
(	596	)	,
(	598	)	,
(	599	)	,
(	600	)	,
(	602	)	,
(	603	)	,
(	605	)	,
(	606	)	,
(	608	)	,
(	609	)	,
(	610	)	,
(	612	)	,
(	613	)	,
(	615	)	,
(	616	)	,
(	618	)	,
(	619	)	,
(	621	)	,
(	622	)	,
(	624	)	,
(	625	)	,
(	627	)	,
(	628	)	,
(	630	)	,
(	631	)	,
(	633	)	,
(	635	)	,
(	636	)	,
(	638	)	,
(	639	)	,
(	641	)	,
(	642	)	,
(	644	)	,
(	646	)	,
(	647	)	,
(	649	)	,
(	650	)	,
(	652	)	,
(	654	)	,
(	655	)	,
(	657	)	,
(	659	)	,
(	660	)	,
(	662	)	,
(	664	)	,
(	665	)	,
(	667	)	,
(	669	)	,
(	670	)	,
(	672	)	,
(	674	)	,
(	675	)	,
(	677	)	,
(	679	)	,
(	681	)	,
(	682	)	,
(	684	)	,
(	686	)	,
(	688	)	,
(	689	)	,
(	691	)	,
(	693	)	,
(	695	)	,
(	697	)	,
(	698	)	,
(	700	)	,
(	702	)	,
(	704	)	,
(	706	)	,
(	708	)	,
(	709	)	,
(	711	)	,
(	713	)	,
(	715	)	,
(	717	)	,
(	719	)	,
(	721	)	,
(	723	)	,
(	724	)	,
(	726	)	,
(	728	)	,
(	730	)	,
(	732	)	,
(	734	)	,
(	736	)	,
(	738	)	,
(	740	)	,
(	742	)	,
(	744	)	,
(	746	)	,
(	748	)	,
(	750	)	,
(	752	)	,
(	754	)	,
(	756	)	,
(	758	)	,
(	760	)	,
(	762	)	,
(	764	)	,
(	766	)	,
(	768	)	,
(	770	)	,
(	772	)	,
(	774	)	,
(	776	)	,
(	779	)	,
(	781	)	,
(	783	)	,
(	785	)	,
(	787	)	,
(	789	)	,
(	791	)	,
(	794	)	,
(	796	)	,
(	798	)	,
(	800	)	,
(	802	)	,
(	804	)	,
(	807	)	,
(	809	)	,
(	811	)	,
(	813	)	,
(	815	)	,
(	818	)	,
(	820	)	,
(	822	)	,
(	824	)	,
(	827	)	,
(	829	)	,
(	831	)	,
(	834	)	,
(	836	)	,
(	838	)	,
(	841	)	,
(	843	)	,
(	845	)	,
(	848	)	,
(	850	)	,
(	852	)	,
(	855	)	,
(	857	)	,
(	859	)	,
(	862	)	,
(	864	)	,
(	867	)	,
(	869	)	,
(	871	)	,
(	874	)	,
(	876	)	,
(	879	)	,
(	881	)	,
(	884	)	,
(	886	)	,
(	889	)	,
(	891	)	,
(	894	)	,
(	896	)	,
(	899	)	,
(	901	)	,
(	904	)	,
(	906	)	,
(	909	)	,
(	911	)	,
(	914	)	,
(	916	)	,
(	919	)	,
(	922	)	,
(	924	)	,
(	927	)	,
(	929	)	,
(	932	)	,
(	935	)	,
(	937	)	,
(	940	)	,
(	943	)	,
(	945	)	,
(	948	)	,
(	951	)	,
(	953	)	,
(	956	)	,
(	959	)	,
(	961	)	,
(	964	)	,
(	967	)	,
(	970	)	,
(	972	)	,
(	975	)	,
(	978	)	,
(	981	)	,
(	983	)	,
(	986	)	,
(	989	)	,
(	992	)	,
(	995	)	,
(	997	)	,
(	1000	)	,
(	1003	)	,
(	1006	)	,
(	1009	)	,
(	1012	)	,
(	1015	)	,
(	1018	)	,
(	1020	)	,
(	1023	)	,
(	1026	)	,
(	1029	)	,
(	1032	)	,
(	1035	)	,
(	1038	)	,
(	1041	)	,
(	1044	)	,
(	1047	)	,
(	1050	)	,
(	1053	)	,
(	1056	)	,
(	1059	)	,
(	1062	)	,
(	1065	)	,
(	1068	)	,
(	1071	)	,
(	1074	)	,
(	1077	)	,
(	1080	)	,
(	1083	)	,
(	1087	)	,
(	1090	)	,
(	1093	)	,
(	1096	)	,
(	1099	)	,
(	1102	)	,
(	1105	)	,
(	1108	)	,
(	1112	)	,
(	1115	)	,
(	1118	)	,
(	1121	)	,
(	1124	)	,
(	1128	)	,
(	1131	)	,
(	1134	)	,
(	1137	)	,
(	1141	)	,
(	1144	)	,
(	1147	)	,
(	1150	)	,
(	1154	)	,
(	1157	)	,
(	1160	)	,
(	1164	)	,
(	1167	)	,
(	1170	)	,
(	1174	)	,
(	1177	)	,
(	1181	)	,
(	1184	)	,
(	1187	)	,
(	1191	)	,
(	1194	)	,
(	1198	)	,
(	1201	)	,
(	1204	)	,
(	1208	)	,
(	1211	)	,
(	1215	)	,
(	1218	)	,
(	1222	)	,
(	1225	)	,
(	1229	)	,
(	1232	)	,
(	1236	)	,
(	1239	)	,
(	1243	)	,
(	1247	)	,
(	1250	)	,
(	1254	)	,
(	1257	)	,
(	1261	)	,
(	1265	)	,
(	1268	)	,
(	1272	)	,
(	1275	)	,
(	1279	)	,
(	1283	)	,
(	1286	)	,
(	1290	)	,
(	1294	)	,
(	1297	)	,
(	1301	)	,
(	1305	)	,
(	1309	)	,
(	1312	)	,
(	1316	)	,
(	1320	)	,
(	1324	)	,
(	1328	)	,
(	1331	)	,
(	1335	)	,
(	1339	)	,
(	1343	)	,
(	1347	)	,
(	1350	)	,
(	1354	)	,
(	1358	)	,
(	1362	)	,
(	1366	)	,
(	1370	)	,
(	1374	)	,
(	1378	)	,
(	1382	)	,
(	1386	)	,
(	1390	)	,
(	1394	)	,
(	1398	)	,
(	1402	)	,
(	1406	)	,
(	1410	)	,
(	1414	)	,
(	1418	)	,
(	1422	)	,
(	1426	)	,
(	1430	)	,
(	1434	)	,
(	1438	)	,
(	1442	)	,
(	1446	)	,
(	1450	)	,
(	1454	)	,
(	1459	)	,
(	1463	)	,
(	1467	)	,
(	1471	)	,
(	1475	)	,
(	1479	)	,
(	1484	)	,
(	1488	)	,
(	1492	)	,
(	1496	)	,
(	1501	)	,
(	1505	)	,
(	1509	)	,
(	1513	)	,
(	1518	)	,
(	1522	)	,
(	1526	)	,
(	1531	)	,
(	1535	)	,
(	1539	)	,
(	1544	)	,
(	1548	)	,
(	1552	)	,
(	1557	)	,
(	1561	)	,
(	1566	)	,
(	1570	)	,
(	1575	)	,
(	1579	)	,
(	1584	)	,
(	1588	)	,
(	1592	)	,
(	1597	)	,
(	1602	)	,
(	1606	)	,
(	1611	)	,
(	1615	)	,
(	1620	)	,
(	1624	)	,
(	1629	)	,
(	1633	)	,
(	1638	)	,
(	1643	)	,
(	1647	)	,
(	1652	)	,
(	1657	)	,
(	1661	)	,
(	1666	)	,
(	1671	)	,
(	1675	)	,
(	1680	)	,
(	1685	)	,
(	1690	)	,
(	1694	)	,
(	1699	)	,
(	1704	)	,
(	1709	)	,
(	1713	)	,
(	1718	)	,
(	1723	)	,
(	1728	)	,
(	1733	)	,
(	1738	)	,
(	1742	)	,
(	1747	)	,
(	1752	)	,
(	1757	)	,
(	1762	)	,
(	1767	)	,
(	1772	)	,
(	1777	)	,
(	1782	)	,
(	1787	)	,
(	1792	)	,
(	1797	)	,
(	1802	)	,
(	1807	)	,
(	1812	)	,
(	1817	)	,
(	1822	)	,
(	1827	)	,
(	1832	)	,
(	1837	)	,
(	1842	)	,
(	1848	)	,
(	1853	)	,
(	1858	)	,
(	1863	)	,
(	1868	)	,
(	1873	)	,
(	1879	)	,
(	1884	)	,
(	1889	)	,
(	1894	)	,
(	1899	)	,
(	1905	)	,
(	1910	)	,
(	1915	)	,
(	1921	)	,
(	1926	)	,
(	1931	)	,
(	1937	)	,
(	1942	)	,
(	1947	)	,
(	1953	)	,
(	1958	)	,
(	1963	)	,
(	1969	)	,
(	1974	)	,
(	1980	)	,
(	1985	)	,
(	1991	)	,
(	1996	)	,
(	2002	)	,
(	2007	)	,
(	2013	)	,
(	2018	)	,
(	2024	)	,
(	2029	)	,
(	2035	)	,
(	2041	)	,
(	2046	)	,
(	2052	)	,
(	2057	)	,
(	2063	)	,
(	2069	)	,
(	2074	)	,
(	2080	)	,
(	2086	)	,
(	2091	)	,
(	2097	)	,
(	2103	)	,
(	2109	)	,
(	2114	)	,
(	2120	)	,
(	2126	)	,
(	2132	)	,
(	2138	)	,
(	2143	)	,
(	2149	)	,
(	2155	)	,
(	2161	)	,
(	2167	)	,
(	2173	)	,
(	2179	)	,
(	2185	)	,
(	2191	)	,
(	2196	)	,
(	2202	)	,
(	2208	)	,
(	2214	)	,
(	2220	)	,
(	2226	)	,
(	2232	)	,
(	2238	)	,
(	2245	)	,
(	2251	)	,
(	2257	)	,
(	2263	)	,
(	2269	)	,
(	2275	)	,
(	2281	)	,
(	2287	)	,
(	2294	)	,
(	2300	)	,
(	2306	)	,
(	2312	)	,
(	2318	)	,
(	2325	)	,
(	2331	)	,
(	2337	)	,
(	2343	)	,
(	2350	)	,
(	2356	)	,
(	2362	)	,
(	2369	)	,
(	2375	)	,
(	2381	)	,
(	2388	)	,
(	2394	)	,
(	2401	)	,
(	2407	)	,
(	2413	)	,
(	2420	)	,
(	2426	)	,
(	2433	)	,
(	2439	)	,
(	2446	)	,
(	2452	)	,
(	2459	)	,
(	2465	)	,
(	2472	)	,
(	2479	)	,
(	2485	)	,
(	2492	)	,
(	2498	)	,
(	2505	)	,
(	2512	)	,
(	2518	)	,
(	2525	)	,
(	2532	)	,
(	2539	)	,
(	2545	)	,
(	2552	)	,
(	2559	)	,
(	2566	)	,
(	2572	)	,
(	2579	)	,
(	2586	)	,
(	2593	)	,
(	2600	)	,
(	2606	)	,
(	2613	)	,
(	2620	)	,
(	2627	)	,
(	2634	)	,
(	2641	)	,
(	2648	)	,
(	2655	)	,
(	2662	)	,
(	2669	)	,
(	2676	)	,
(	2683	)	,
(	2690	)	,
(	2697	)	,
(	2704	)	,
(	2711	)	,
(	2718	)	,
(	2725	)	,
(	2733	)	,
(	2740	)	,
(	2747	)	,
(	2754	)	,
(	2761	)	,
(	2769	)	,
(	2776	)	,
(	2783	)	,
(	2790	)	,
(	2798	)	,
(	2805	)	,
(	2812	)	,
(	2819	)	,
(	2827	)	,
(	2834	)	,
(	2841	)	,
(	2849	)	,
(	2856	)	,
(	2864	)	,
(	2871	)	,
(	2879	)	,
(	2886	)	,
(	2893	)	,
(	2901	)	,
(	2908	)	,
(	2916	)	,
(	2924	)	,
(	2931	)	,
(	2939	)	,
(	2946	)	,
(	2954	)	,
(	2961	)	,
(	2969	)	,
(	2977	)	,
(	2984	)	,
(	2992	)	,
(	3000	)	,
(	3007	)	,
(	3015	)	,
(	3023	)	,
(	3031	)	,
(	3038	)	,
(	3046	)	,
(	3054	)	,
(	3062	)	,
(	3070	)	,
(	3078	)	,
(	3085	)	,
(	3093	)	,
(	3101	)	,
(	3109	)	,
(	3117	)	,
(	3125	)	,
(	3133	)	,
(	3141	)	,
(	3149	)	,
(	3157	)	,
(	3165	)	,
(	3173	)	,
(	3181	)	,
(	3189	)	,
(	3197	)	,
(	3206	)	,
(	3214	)	,
(	3222	)	,
(	3230	)	,
(	3238	)	,
(	3246	)	,
(	3255	)	,
(	3263	)	,
(	3271	)	,
(	3279	)	,
(	3288	)	,
(	3296	)	,
(	3304	)	,
(	3313	)	,
(	3321	)	,
(	3329	)	,
(	3338	)	,
(	3346	)	,
(	3355	)	,
(	3363	)	,
(	3371	)	,
(	3380	)	,
(	3388	)	,
(	3397	)	,
(	3405	)	,
(	3414	)	,
(	3423	)	,
(	3431	)	,
(	3440	)	,
(	3448	)	,
(	3457	)	,
(	3466	)	,
(	3474	)	,
(	3483	)	,
(	3492	)	,
(	3500	)	,
(	3509	)	,
(	3518	)	,
(	3527	)	,
(	3535	)	,
(	3544	)	,
(	3553	)	,
(	3562	)	,
(	3571	)	,
(	3580	)	,
(	3588	)	,
(	3597	)	,
(	3606	)	,
(	3615	)	,
(	3624	)	,
(	3633	)	,
(	3642	)	,
(	3651	)	,
(	3660	)	,
(	3669	)	,
(	3678	)	,
(	3687	)	,
(	3696	)	,
(	3706	)	,
(	3715	)	,
(	3724	)	,
(	3733	)	,
(	3742	)	,
(	3751	)	,
(	3761	)	,
(	3770	)	,
(	3779	)	,
(	3788	)	,
(	3798	)	,
(	3807	)	,
(	3816	)	,
(	3826	)	,
(	3835	)	,
(	3844	)	,
(	3854	)	,
(	3863	)	,
(	3873	)	,
(	3882	)	,
(	3892	)	,
(	3901	)	,
(	3911	)	,
(	3920	)	,
(	3930	)	,
(	3939	)	,
(	3949	)	,
(	3958	)	,
(	3968	)	,
(	3978	)	,
(	3987	)	,
(	3997	)	,
(	4007	)	,
(	4016	)	,
(	4026	)	,
(	4036	)	,
(	4046	)	,
(	4055	)	,
(	4065	)	,
(	4075	)	,
(	4085	)	,
(	4095	)	,
(	4105	)	,
(	4115	)	,
(	4124	)	,
(	4134	)	,
(	4144	)	,
(	4154	)	,
(	4164	)	,
(	4174	)	,
(	4184	)	,
(	4194	)	,
(	4204	)	,
(	4215	)	,
(	4225	)	,
(	4235	)	,
(	4245	)	,
(	4255	)	,
(	4265	)	,
(	4276	)	,
(	4286	)	,
(	4296	)	,
(	4306	)	,
(	4317	)	,
(	4327	)	,
(	4337	)	,
(	4347	)	,
(	4358	)	,
(	4368	)	,
(	4379	)	,
(	4389	)	,
(	4399	)	,
(	4410	)	,
(	4420	)	,
(	4431	)	,
(	4441	)	,
(	4452	)	,
(	4462	)	,
(	4473	)	,
(	4484	)	,
(	4494	)	,
(	4505	)	,
(	4515	)	,
(	4526	)	,
(	4537	)	,
(	4548	)	,
(	4558	)	,
(	4569	)	,
(	4580	)	,
(	4591	)	,
(	4601	)	,
(	4612	)	,
(	4623	)	,
(	4634	)	,
(	4645	)	,
(	4656	)	,
(	4667	)	,
(	4678	)	,
(	4688	)	,
(	4699	)	,
(	4710	)	,
(	4721	)	,
(	4733	)	,
(	4744	)	,
(	4755	)	,
(	4766	)	,
(	4777	)	,
(	4788	)	,
(	4799	)	,
(	4810	)	,
(	4822	)	,
(	4833	)	,
(	4844	)	,
(	4855	)	,
(	4867	)	,
(	4878	)	,
(	4889	)	,
(	4901	)	,
(	4912	)	,
(	4923	)	,
(	4935	)	,
(	4946	)	,
(	4958	)	,
(	4969	)	,
(	4981	)	,
(	4992	)	,
(	5004	)	,
(	5015	)	,
(	5027	)	,
(	5038	)	,
(	5050	)	,
(	5062	)	,
(	5073	)	,
(	5085	)	,
(	5097	)	,
(	5108	)	,
(	5120	)	,
(	5132	)	,
(	5144	)	,
(	5155	)	,
(	5167	)	,
(	5179	)	,
(	5191	)	,
(	5203	)	,
(	5215	)	,
(	5227	)	,
(	5239	)	,
(	5251	)	,
(	5263	)	,
(	5275	)	,
(	5287	)	,
(	5299	)	,
(	5311	)	,
(	5323	)	,
(	5335	)	,
(	5347	)	,
(	5359	)	,
(	5371	)	,
(	5384	)	,
(	5396	)	,
(	5408	)	,
(	5420	)	,
(	5433	)	,
(	5445	)	,
(	5457	)	,
(	5470	)	,
(	5482	)	,
(	5494	)	,
(	5507	)	,
(	5519	)	,
(	5532	)	,
(	5544	)	,
(	5557	)	,
(	5569	)	,
(	5582	)	,
(	5594	)	,
(	5607	)	,
(	5620	)	,
(	5632	)	,
(	5645	)	,
(	5658	)	,
(	5670	)	,
(	5683	)	,
(	5696	)	,
(	5709	)	,
(	5721	)	,
(	5734	)	,
(	5747	)	,
(	5760	)	,
(	5773	)	,
(	5786	)	,
(	5799	)	,
(	5812	)	,
(	5824	)	,
(	5837	)	,
(	5850	)	,
(	5864	)	,
(	5877	)	,
(	5890	)	,
(	5903	)	,
(	5916	)	,
(	5929	)	,
(	5942	)	,
(	5955	)	,
(	5969	)	,
(	5982	)	,
(	5995	)	,
(	6008	)	,
(	6022	)	,
(	6035	)	,
(	6048	)	,
(	6062	)	,
(	6075	)	,
(	6089	)	,
(	6102	)	,
(	6115	)	,
(	6129	)	,
(	6142	)	,
(	6156	)	,
(	6170	)	,
(	6183	)	,
(	6197	)	,
(	6210	)	,
(	6224	)	,
(	6238	)	,
(	6251	)	,
(	6265	)	,
(	6279	)	,
(	6293	)	,
(	6306	)	,
(	6320	)	,
(	6334	)	,
(	6348	)	,
(	6362	)	,
(	6376	)	,
(	6389	)	,
(	6403	)	,
(	6417	)	,
(	6431	)	,
(	6445	)	,
(	6459	)	,
(	6474	)	,
(	6488	)	,
(	6502	)	,
(	6516	)	,
(	6530	)	,
(	6544	)	,
(	6558	)	,
(	6573	)	,
(	6587	)	,
(	6601	)	,
(	6615	)	,
(	6630	)	,
(	6644	)	,
(	6658	)	,
(	6673	)	,
(	6687	)	,
(	6702	)	,
(	6716	)	,
(	6731	)	,
(	6745	)	,
(	6760	)	,
(	6774	)	,
(	6789	)	,
(	6803	)	,
(	6818	)	,
(	6833	)	,
(	6847	)	,
(	6862	)	,
(	6877	)	,
(	6892	)	,
(	6906	)	,
(	6921	)	,
(	6936	)	,
(	6951	)	,
(	6966	)	,
(	6981	)	,
(	6996	)	,
(	7010	)	,
(	7025	)	,
(	7040	)	,
(	7055	)	,
(	7071	)	,
(	7086	)	,
(	7101	)	,
(	7116	)	,
(	7131	)	,
(	7146	)	,
(	7161	)	,
(	7176	)	,
(	7192	)	,
(	7207	)	,
(	7222	)	,
(	7238	)	,
(	7253	)	,
(	7268	)	,
(	7284	)	,
(	7299	)	,
(	7315	)	,
(	7330	)	,
(	7345	)	,
(	7361	)	,
(	7377	)	,
(	7392	)	,
(	7408	)	,
(	7423	)	,
(	7439	)	,
(	7455	)	,
(	7470	)	,
(	7486	)	,
(	7502	)	,
(	7518	)	,
(	7533	)	,
(	7549	)	,
(	7565	)	,
(	7581	)	,
(	7597	)	,
(	7613	)	,
(	7629	)	,
(	7645	)	,
(	7661	)	,
(	7677	)	,
(	7693	)	,
(	7709	)	,
(	7725	)	,
(	7741	)	,
(	7757	)	,
(	7773	)	,
(	7789	)	,
(	7806	)	,
(	7822	)	,
(	7838	)	,
(	7854	)	,
(	7871	)	,
(	7887	)	,
(	7903	)	,
(	7920	)	,
(	7936	)	,
(	7953	)	,
(	7969	)	,
(	7986	)	,
(	8002	)	,
(	8019	)	,
(	8035	)	,
(	8052	)	,
(	8069	)	,
(	8085	)	,
(	8102	)	,
(	8119	)	,
(	8135	)	,
(	8152	)	,
(	8169	)	,
(	8186	)	,
(	8203	)	,
(	8219	)	,
(	8236	)	,
(	8253	)	,
(	8270	)	,
(	8287	)	,
(	8304	)	,
(	8321	)	,
(	8338	)	,
(	8355	)	,
(	8373	)	,
(	8390	)	,
(	8407	)	,
(	8424	)	,
(	8441	)	,
(	8458	)	,
(	8476	)	,
(	8493	)	,
(	8510	)	,
(	8528	)	,
(	8545	)	,
(	8562	)	,
(	8580	)	,
(	8597	)	,
(	8615	)	,
(	8632	)	,
(	8650	)	,
(	8667	)	,
(	8685	)	,
(	8703	)	,
(	8720	)	,
(	8738	)	,
(	8756	)	,
(	8773	)	,
(	8791	)	,
(	8809	)	,
(	8827	)	,
(	8845	)	,
(	8862	)	,
(	8880	)	,
(	8898	)	,
(	8916	)	,
(	8934	)	,
(	8952	)	,
(	8970	)	,
(	8988	)	,
(	9006	)	,
(	9024	)	,
(	9043	)	,
(	9061	)	,
(	9079	)	,
(	9097	)	,
(	9115	)	,
(	9134	)	,
(	9152	)	,
(	9170	)	,
(	9189	)	,
(	9207	)	,
(	9225	)	,
(	9244	)	,
(	9262	)	,
(	9281	)	,
(	9299	)	,
(	9318	)	,
(	9337	)	,
(	9355	)	,
(	9374	)	,
(	9392	)	,
(	9411	)	,
(	9430	)	,
(	9449	)	,
(	9467	)	,
(	9486	)	,
(	9505	)	,
(	9524	)	,
(	9543	)	,
(	9562	)	,
(	9581	)	,
(	9600	)	,
(	9619	)	,
(	9638	)	,
(	9657	)	,
(	9676	)	,
(	9695	)	,
(	9714	)	,
(	9733	)	,
(	9752	)	,
(	9772	)	,
(	9791	)	,
(	9810	)	,
(	9830	)	,
(	9849	)	,
(	9868	)	,
(	9888	)	,
(	9907	)	,
(	9927	)	,
(	9946	)	,
(	9966	)	,
(	9985	)	,
(	10005	)	,
(	10024	)	,
(	10044	)	,
(	10064	)	,
(	10083	)	,
(	10103	)	,
(	10123	)	,
(	10143	)	,
(	10162	)	,
(	10182	)	,
(	10202	)	,
(	10222	)	,
(	10242	)	,
(	10262	)	,
(	10282	)	,
(	10302	)	,
(	10322	)	,
(	10342	)	,
(	10362	)	,
(	10382	)	,
(	10402	)	,
(	10423	)	,
(	10443	)	,
(	10463	)	,
(	10483	)	,
(	10504	)	,
(	10524	)	,
(	10544	)	,
(	10565	)	,
(	10585	)	,
(	10606	)	,
(	10626	)	,
(	10647	)	,
(	10667	)	,
(	10688	)	,
(	10708	)	,
(	10729	)	,
(	10750	)	,
(	10770	)	,
(	10791	)	,
(	10812	)	,
(	10833	)	,
(	10854	)	,
(	10874	)	,
(	10895	)	,
(	10916	)	,
(	10937	)	,
(	10958	)	,
(	10979	)	,
(	11000	)	,
(	11021	)	,
(	11042	)	,
(	11063	)	,
(	11085	)	,
(	11106	)	,
(	11127	)	,
(	11148	)	,
(	11170	)	,
(	11191	)	,
(	11212	)	,
(	11234	)	,
(	11255	)	,
(	11276	)	,
(	11298	)	,
(	11319	)	,
(	11341	)	,
(	11362	)	,
(	11384	)	,
(	11406	)	,
(	11427	)	,
(	11449	)	,
(	11471	)	,
(	11492	)	,
(	11514	)	,
(	11536	)	,
(	11558	)	,
(	11580	)	,
(	11602	)	,
(	11623	)	,
(	11645	)	,
(	11667	)	,
(	11689	)	,
(	11711	)	,
(	11734	)	,
(	11756	)	,
(	11778	)	,
(	11800	)	,
(	11822	)	,
(	11844	)	,
(	11867	)	,
(	11889	)	,
(	11911	)	,
(	11934	)	,
(	11956	)	,
(	11979	)	,
(	12001	)	,
(	12023	)	,
(	12046	)	,
(	12069	)	,
(	12091	)	,
(	12114	)	,
(	12136	)	,
(	12159	)	,
(	12182	)	,
(	12205	)	,
(	12227	)	,
(	12250	)	,
(	12273	)	,
(	12296	)	,
(	12319	)	,
(	12342	)	,
(	12365	)	,
(	12388	)	,
(	12411	)	,
(	12434	)	,
(	12457	)	,
(	12480	)	,
(	12503	)	,
(	12526	)	,
(	12550	)	,
(	12573	)	,
(	12596	)	,
(	12619	)	,
(	12643	)	,
(	12666	)	,
(	12690	)	,
(	12713	)	,
(	12737	)	,
(	12760	)	,
(	12784	)	,
(	12807	)	,
(	12831	)	,
(	12854	)	,
(	12878	)	,
(	12902	)	,
(	12926	)	,
(	12949	)	,
(	12973	)	,
(	12997	)	,
(	13021	)	,
(	13045	)	,
(	13069	)	,
(	13093	)	,
(	13117	)	,
(	13141	)	,
(	13165	)	,
(	13189	)	,
(	13213	)	,
(	13237	)	,
(	13262	)	,
(	13286	)	,
(	13310	)	,
(	13334	)	,
(	13359	)	,
(	13383	)	,
(	13408	)	,
(	13432	)	,
(	13457	)	,
(	13481	)	,
(	13506	)	,
(	13530	)	,
(	13555	)	,
(	13579	)	,
(	13604	)	,
(	13629	)	,
(	13654	)	,
(	13678	)	,
(	13703	)	,
(	13728	)	,
(	13753	)	,
(	13778	)	,
(	13803	)	,
(	13828	)	,
(	13853	)	,
(	13878	)	,
(	13903	)	,
(	13928	)	,
(	13953	)	,
(	13978	)	,
(	14004	)	,
(	14029	)	,
(	14054	)	,
(	14079	)	,
(	14105	)	,
(	14130	)	,
(	14156	)	,
(	14181	)	,
(	14207	)	,
(	14232	)	,
(	14258	)	,
(	14283	)	,
(	14309	)	,
(	14335	)	,
(	14360	)	,
(	14386	)	,
(	14412	)	,
(	14438	)	,
(	14464	)	,
(	14489	)	,
(	14515	)	,
(	14541	)	,
(	14567	)	,
(	14593	)	,
(	14619	)	,
(	14645	)	,
(	14672	)	,
(	14698	)	,
(	14724	)	,
(	14750	)	,
(	14776	)	,
(	14803	)	,
(	14829	)	,
(	14855	)	,
(	14882	)	,
(	14908	)	,
(	14935	)	,
(	14961	)	,
(	14988	)	,
(	15014	)	,
(	15041	)	,
(	15068	)	,
(	15094	)	,
(	15121	)	,
(	15148	)	,
(	15175	)	,
(	15201	)	,
(	15228	)	,
(	15255	)	,
(	15282	)	,
(	15309	)	,
(	15336	)	,
(	15363	)	,
(	15390	)	,
(	15417	)	,
(	15444	)	,
(	15472	)	,
(	15499	)	,
(	15526	)	,
(	15553	)	,
(	15581	)	,
(	15608	)	,
(	15635	)	,
(	15663	)	,
(	15690	)	,
(	15718	)	,
(	15745	)	,
(	15773	)	,
(	15801	)	,
(	15828	)	,
(	15856	)	,
(	15884	)	,
(	15911	)	,
(	15939	)	,
(	15967	)	,
(	15995	)	,
(	16023	)	,
(	16051	)	,
(	16079	)	,
(	16107	)	,
(	16135	)	,
(	16163	)	,
(	16191	)	,
(	16219	)	,
(	16247	)	,
(	16276	)	,
(	16304	)	,
(	16332	)	,
(	16361	)	,
(	16389	)	,
(	16417	)	,
(	16446	)	,
(	16474	)	,
(	16503	)	,
(	16532	)	,
(	16560	)	,
(	16589	)	,
(	16617	)	,
(	16646	)	,
(	16675	)	,
(	16704	)	,
(	16733	)	,
(	16761	)	,
(	16790	)	,
(	16819	)	,
(	16848	)	,
(	16877	)

);


end package LUT_pkg;
